.SUBCKT MAC in1_IFM[3] in1_IFM[2] in1_IFM[1] in1_IFM[0] in2_IFM[3] in2_IFM[2] in2_IFM[1] in2_IFM[0] out[9] out[8] out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0] clk rst_n in_valid out_valid
Xcstate_reg_0_ n108 clk n238 n138 n106 ASYNC_DFFHx1_ASAP7_75t_R
Xcstate_reg_1_ n107 clk n238 n128 n105 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_3_ N25 clk n238 n167 n104 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_2_ N24 clk n238 n148 n103 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_1_ N23 clk n238 n125 n102 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_0_ N22 clk n238 n119 n101 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_3_ N21 clk n238 n124 n100 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_2_ N20 clk n238 n121 n99 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_1_ N19 clk n238 n116 n98 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_0_ N18 clk n238 n156 n97 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_7_ add_x_7_n6 clk n238 n145 n96 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_6_ add_x_8_n6 clk n238 n137 n95 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_5_ add_x_9_n6 clk n238 n154 n94 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_4_ add_x_10_n6 clk n238 n146 n93 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_3_ add_x_11_n6 clk n238 n142 n92 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_2_ add_x_12_n6 clk n238 n122 n91 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_1_ add_x_6_n6 clk n238 n141 n90 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_0_ fprod_0_ clk n238 n131 n89 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_8_ temp_1 clk n238 n117 n88 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_7_ temp_0[7] clk n238 n129 n87 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_6_ temp_0[6] clk n238 n140 n86 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_5_ temp_0[5] clk n238 n157 n85 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_4_ temp_0[4] clk n238 n127 n84 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_3_ temp_0[3] clk n238 n126 n83 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_2_ temp_0[2] clk n238 n155 n82 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_1_ temp_0[1] clk n238 n115 n81 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_0_ temp_0[0] clk n238 n166 n80 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_8_ N37 clk n238 n130 n79 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_7_ N36 clk n238 n151 n78 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_6_ N35 clk n238 n123 n77 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_5_ N34 clk n238 n118 n76 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_4_ N33 clk n238 n120 n75 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_3_ N32 clk n238 n147 n74 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_2_ N31 clk n238 n144 n73 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_1_ N30 clk n238 n132 n72 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_0_ N29 clk n238 n139 n71 ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg n218 clk n238 n109 n69 ASYNC_DFFHx1_ASAP7_75t_R
XU128 n143 n226 add_x_9_n6 NOR2xp33_ASAP7_75t_R
XU129 in_valid in2_IFM[1] N23 AND2x2_ASAP7_75t_R
XU130 in_valid in2_IFM[2] N24 AND2x2_ASAP7_75t_R
XU131 in_valid in2_IFM[0] N22 AND2x2_ASAP7_75t_R
XU132 in_valid in2_IFM[3] N25 AND2x2_ASAP7_75t_R
XU133 in_valid in1_IFM[2] N20 AND2x2_ASAP7_75t_R
XU134 in_valid in1_IFM[1] N19 AND2x2_ASAP7_75t_R
XU135 in_valid in1_IFM[0] N18 AND2x2_ASAP7_75t_R
XU136 n235 n162 INVx3_ASAP7_75t_R
XU137 n158 n236 INVx3_ASAP7_75t_R
XU138 n195 n194 n223 NOR2xp33_ASAP7_75t_R
XU139 n134 n183 n188 NOR2xp33_ASAP7_75t_R
XU140 n104 n99 n189 NOR2xp33_ASAP7_75t_R
XU141 n100 n103 n190 NOR2xp33_ASAP7_75t_R
XU142 n181 n180 n159 XOR2xp5_ASAP7_75t_R
XU143 n173 n172 n191 NOR2xp33_ASAP7_75t_R
XU144 n111 TIEHIx1_ASAP7_75t_R
XU145 n111 out[9] INVx1_ASAP7_75t_R
XU146 n218 n112 INVx4_ASAP7_75t_R
XU147 n162 n236 n218 AND2x6_ASAP7_75t_R
XU148 n105 n235 BUFx5_ASAP7_75t_R
XU149 n106 n158 BUFx5_ASAP7_75t_R
XU150 n186 n185 n187 NOR2xp33_ASAP7_75t_R
XU151 n103 n98 n177 NOR2xp33_ASAP7_75t_R
XU152 n202 n201 n227 NOR2xp33_ASAP7_75t_R
XU153 in_valid in1_IFM[3] N21 AND2x2_ASAP7_75t_R
XU154 n150 n203 add_x_7_n6 NAND2xp5_ASAP7_75t_R
XU155 n233 n219 n221 NAND2xp5_ASAP7_75t_R
XU156 n152 n207 INVx2_ASAP7_75t_R
XU157 n190 n189 n161 NAND2xp5_ASAP7_75t_R
XU158 n149 n215 INVx2_ASAP7_75t_R
XU159 n153 n211 INVx2_ASAP7_75t_R
XU160 n181 n180 n160 XNOR2xp5_ASAP7_75t_R
XU161 n188 n187 n199 XNOR2xp5_ASAP7_75t_R
XU162 n179 n184 n113 XOR2xp5_ASAP7_75t_R
XU163 n179 n184 n197 XNOR2xp5_ASAP7_75t_R
XU164 n225 n224 n114 NAND2xp33_ASAP7_75t_R
XU165 rst_n n115 INVx8_ASAP7_75t_R
XU166 rst_n n116 INVx8_ASAP7_75t_R
XU167 rst_n n117 INVx8_ASAP7_75t_R
XU168 rst_n n118 INVx8_ASAP7_75t_R
XU169 rst_n n119 INVx8_ASAP7_75t_R
XU170 rst_n n120 INVx8_ASAP7_75t_R
XU171 rst_n n121 INVx8_ASAP7_75t_R
XU172 rst_n n122 INVx8_ASAP7_75t_R
XU173 rst_n n123 INVx8_ASAP7_75t_R
XU174 rst_n n124 INVx8_ASAP7_75t_R
XU175 rst_n n125 INVx8_ASAP7_75t_R
XU176 rst_n n126 INVx8_ASAP7_75t_R
XU177 rst_n n127 INVx8_ASAP7_75t_R
XU178 rst_n n128 INVx8_ASAP7_75t_R
XU179 rst_n n129 INVx8_ASAP7_75t_R
XU180 rst_n n130 INVx8_ASAP7_75t_R
XU181 rst_n n131 INVx8_ASAP7_75t_R
XU182 rst_n n132 INVx8_ASAP7_75t_R
XU183 n188 n187 n133 XOR2xp5_ASAP7_75t_R
XU184 n221 n220 n134 NOR2xp33_ASAP7_75t_R
XU185 n182 n159 n135 XOR2xp5_ASAP7_75t_R
XU186 n225 n224 n143 AND2x2_ASAP7_75t_R
XU187 n190 n189 n136 AND2x2_ASAP7_75t_R
XU188 rst_n n137 INVx8_ASAP7_75t_R
XU189 rst_n n138 INVx8_ASAP7_75t_R
XU190 rst_n n139 INVx8_ASAP7_75t_R
XU191 rst_n n140 INVx8_ASAP7_75t_R
XU192 rst_n n141 INVx8_ASAP7_75t_R
XU193 rst_n n142 INVx8_ASAP7_75t_R
XU194 n188 n161 n150 OR2x2_ASAP7_75t_R
XU195 rst_n n144 INVx8_ASAP7_75t_R
XU196 rst_n n145 INVx8_ASAP7_75t_R
XU197 n221 n220 n184 OR2x2_ASAP7_75t_R
XU198 n182 n159 n196 XNOR2xp5_ASAP7_75t_R
XU199 rst_n n146 INVx8_ASAP7_75t_R
XU200 rst_n n147 INVx8_ASAP7_75t_R
XU201 rst_n n148 INVx8_ASAP7_75t_R
XU202 n95 n149 BUFx5_ASAP7_75t_R
XU203 rst_n n151 INVx8_ASAP7_75t_R
XU204 n91 n152 BUFx5_ASAP7_75t_R
XU205 n93 n153 BUFx5_ASAP7_75t_R
XU206 rst_n n154 INVx8_ASAP7_75t_R
XU207 rst_n n155 INVx8_ASAP7_75t_R
XU208 rst_n n156 INVx8_ASAP7_75t_R
XU209 rst_n n157 INVx8_ASAP7_75t_R
XU210 n86 n214 BUFx5_ASAP7_75t_R
XU211 n214 n163 INVx4_ASAP7_75t_R
XU212 n84 n210 BUFx5_ASAP7_75t_R
XU213 n210 n164 INVx4_ASAP7_75t_R
XU214 n82 n206 BUFx5_ASAP7_75t_R
XU215 n206 n165 INVx4_ASAP7_75t_R
XU216 rst_n n166 INVx8_ASAP7_75t_R
XU217 rst_n n167 INVx8_ASAP7_75t_R
XU218 rst_n n109 INVx8_ASAP7_75t_R
XU219 n238 TIELOx1_ASAP7_75t_R
XU220 n102 n98 n97 n101 n233 NOR4xp25_ASAP7_75t_R
XU221 n103 n97 n170 NOR2xp33_ASAP7_75t_R
XU222 n102 n98 n169 NOR2xp33_ASAP7_75t_R
XU223 n99 n101 n168 NOR2xp33_ASAP7_75t_R
XU224 n169 n168 n171 HAxp5_ASAP7_75t_R
XU225 n170 n171 n219 HAxp5_ASAP7_75t_R
XU226 n99 n102 n98 n101 n173 NOR4xp25_ASAP7_75t_R
XU227 n103 n97 n171 n172 NOR3xp33_ASAP7_75t_R
XU228 n104 n97 n174 NOR2xp33_ASAP7_75t_R
XU229 n191 n174 n193 HAxp5_ASAP7_75t_R
XU230 n99 n102 n178 NOR2xp33_ASAP7_75t_R
XU231 n100 n101 n176 NOR2xp33_ASAP7_75t_R
XU232 n178 n176 n175 HAxp5_ASAP7_75t_R
XU233 n177 n175 n192 HAxp5_ASAP7_75t_R
XU234 n193 n192 n220 HAxp5_ASAP7_75t_R
XU235 n178 n177 n176 n179 MAJIxp5_ASAP7_75t_R
XU236 n104 n98 n182 NOR2xp33_ASAP7_75t_R
XU237 n103 n99 n181 NOR2xp33_ASAP7_75t_R
XU238 n100 n102 n180 NOR2xp33_ASAP7_75t_R
XU239 n197 n196 n183 NOR2xp33_ASAP7_75t_R
XU240 n188 n161 n202 NOR2xp33_ASAP7_75t_R
XU241 n100 n104 n228 NOR2xp33_ASAP7_75t_R
XU242 n100 n103 n99 n102 n186 NOR4xp25_ASAP7_75t_R
XU243 n104 n98 n160 n185 NOR3xp33_ASAP7_75t_R
XU244 n190 n189 n198 HAxp5_ASAP7_75t_R
XU245 n198 n133 n225 HAxp5_ASAP7_75t_R
XU246 n104 n97 n191 n195 NOR3xp33_ASAP7_75t_R
XU247 n193 n192 n194 AND2x2_ASAP7_75t_R
XU248 n135 n113 n222 HAxp5_ASAP7_75t_R
XU249 n223 n222 n224 NOR2xp33_ASAP7_75t_R
XU250 n199 n198 n200 NOR2xp33_ASAP7_75t_R
XU251 n136 n200 n201 NOR2xp33_ASAP7_75t_R
XU252 n143 n228 n227 n203 MAJIxp5_ASAP7_75t_R
XU253 n69 out_valid INVxp33_ASAP7_75t_R
XU254 n71 out[0] INVxp33_ASAP7_75t_R
XU255 n73 out[2] INVxp33_ASAP7_75t_R
XU256 n74 out[3] INVxp33_ASAP7_75t_R
XU257 n75 out[4] INVxp33_ASAP7_75t_R
XU258 n76 out[5] INVxp33_ASAP7_75t_R
XU259 n77 out[6] INVxp33_ASAP7_75t_R
XU260 n78 out[7] INVxp33_ASAP7_75t_R
XU261 n79 out[8] INVxp33_ASAP7_75t_R
XU262 n72 out[1] INVxp33_ASAP7_75t_R
XU263 n80 n89 temp_0[0] XOR2xp5_ASAP7_75t_R
XU264 n80 n89 n204 OR2x2_ASAP7_75t_R
XU265 n81 n90 n204 temp_0[1] FAx1_ASAP7_75t_R
XU266 n90 n81 n204 n205 MAJIxp5_ASAP7_75t_R
XU267 n152 n205 n165 temp_0[2] FAx1_ASAP7_75t_R
XU268 n207 n205 n165 n208 MAJIxp5_ASAP7_75t_R
XU269 n92 n83 n208 temp_0[3] FAx1_ASAP7_75t_R
XU270 n92 n83 n208 n209 MAJIxp5_ASAP7_75t_R
XU271 n153 n209 n164 temp_0[4] FAx1_ASAP7_75t_R
XU272 n211 n209 n164 n212 MAJIxp5_ASAP7_75t_R
XU273 n94 n85 n212 temp_0[5] FAx1_ASAP7_75t_R
XU274 n94 n85 n212 n213 MAJIxp5_ASAP7_75t_R
XU275 n149 n213 n163 temp_0[6] FAx1_ASAP7_75t_R
XU276 n215 n213 n163 n216 MAJIxp5_ASAP7_75t_R
XU277 n87 n216 n96 temp_0[7] FAx1_ASAP7_75t_R
XU278 n87 n216 n96 n217 MAJIxp5_ASAP7_75t_R
XU279 n88 n217 temp_1 HAxp5_ASAP7_75t_R
XU280 n97 n101 fprod_0_ NOR2xp33_ASAP7_75t_R
XU281 n112 n80 N29 NOR2xp33_ASAP7_75t_R
XU282 n112 n81 N30 NOR2xp33_ASAP7_75t_R
XU283 n206 n112 N31 NOR2xp33_ASAP7_75t_R
XU284 n112 n83 N32 NOR2xp33_ASAP7_75t_R
XU285 n210 n112 N33 NOR2xp33_ASAP7_75t_R
XU286 n112 n85 N34 NOR2xp33_ASAP7_75t_R
XU287 n214 n112 N35 NOR2xp33_ASAP7_75t_R
XU288 n112 n87 N36 NOR2xp33_ASAP7_75t_R
XU289 n112 n88 N37 NOR2xp33_ASAP7_75t_R
XU290 n233 n219 add_x_12_n6 XOR2xp5_ASAP7_75t_R
XU291 n221 n220 add_x_11_n6 XOR2xp5_ASAP7_75t_R
XU292 n223 n222 add_x_10_n6 XOR2xp5_ASAP7_75t_R
XU293 n225 n224 n226 NOR2xp33_ASAP7_75t_R
XU294 n228 n227 n229 XOR2xp5_ASAP7_75t_R
XU295 n229 n114 add_x_8_n6 HAxp5_ASAP7_75t_R
XU296 n98 n101 n231 NOR2xp33_ASAP7_75t_R
XU297 n102 n97 n230 NOR2xp33_ASAP7_75t_R
XU298 n231 n230 n232 NOR2xp33_ASAP7_75t_R
XU299 n233 n232 add_x_6_n6 NOR2xp33_ASAP7_75t_R
XU300 n162 in_valid n234 NOR2xp33_ASAP7_75t_R
XU301 n236 n234 n108 NOR2xp33_ASAP7_75t_R
XU302 n236 n162 n237 NOR2xp33_ASAP7_75t_R
XU303 n218 n237 n107 NOR2xp33_ASAP7_75t_R
.ENDS


