.SUBCKT MAC_v2 VSS VDD  in1_IFM[3] in1_IFM[2] in1_IFM[1] in1_IFM[0] in2_IFM[3] in2_IFM[2] in2_IFM[1] in2_IFM[0] out[9] out[8] out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0] clk rst_n in_valid out_valid
Xcstate_reg_0_ VSS VDD  n42 clk n141 n60 n40 ASYNC_DFFHx1_ASAP7_75t_R
Xcstate_reg_1_ VSS VDD  n41 clk n141 n65 n39 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_3_ VSS VDD  NC25 clk n141 n78 n38 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_2_ VSS VDD  NC24 clk n141 n73 n37 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_1_ VSS VDD  NC23 clk n141 n61 n36 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_0_ VSS VDD  NC22 clk n141 n58 n35 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_3_ VSS VDD  NC21 clk n141 n85 n34 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_2_ VSS VDD  NC20 clk n141 n53 n33 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_1_ VSS VDD  NC19 clk n141 n56 n32 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_0_ VSS VDD  NC18 clk n141 n69 n31 ASYNC_DFFHx1_ASAP7_75t_R
Xtttemp_reg_7_ VSS VDD  NC43 clk n141 n72 n30 ASYNC_DFFHx1_ASAP7_75t_R
Xtttemp_reg_6_ VSS VDD  NC42 clk n141 n84 n29 ASYNC_DFFHx1_ASAP7_75t_R
Xtttemp_reg_5_ VSS VDD  NC41 clk n141 n66 n28 ASYNC_DFFHx1_ASAP7_75t_R
Xtttemp_reg_4_ VSS VDD  NC40 clk n141 n63 n27 ASYNC_DFFHx1_ASAP7_75t_R
Xtttemp_reg_3_ VSS VDD  NC39 clk n141 n67 n26 ASYNC_DFFHx1_ASAP7_75t_R
Xtttemp_reg_2_ VSS VDD  NC38 clk n141 n70 n25 ASYNC_DFFHx1_ASAP7_75t_R
Xtttemp_reg_1_ VSS VDD  NC37 clk n141 n96 n24 ASYNC_DFFHx1_ASAP7_75t_R
Xtttemp_reg_0_ VSS VDD  NC36 clk n141 n80 n23 ASYNC_DFFHx1_ASAP7_75t_R
Xtemp_reg_7_ VSS VDD  NC35 clk n141 n83 n22 ASYNC_DFFHx1_ASAP7_75t_R
Xtemp_reg_6_ VSS VDD  NC34 clk n141 n71 n21 ASYNC_DFFHx1_ASAP7_75t_R
Xtemp_reg_5_ VSS VDD  NC33 clk n141 n75 n20 ASYNC_DFFHx1_ASAP7_75t_R
Xtemp_reg_4_ VSS VDD  NC32 clk n141 n57 n19 ASYNC_DFFHx1_ASAP7_75t_R
Xtemp_reg_3_ VSS VDD  NC31 clk n141 n97 n18 ASYNC_DFFHx1_ASAP7_75t_R
Xtemp_reg_2_ VSS VDD  NC30 clk n141 n62 n17 ASYNC_DFFHx1_ASAP7_75t_R
Xtemp_reg_1_ VSS VDD  NC29 clk n141 n52 n16 ASYNC_DFFHx1_ASAP7_75t_R
Xtemp_reg_0_ VSS VDD  NC28 clk n141 n49 n15 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_7_ VSS VDD  NC52 clk n141 n59 n14 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_6_ VSS VDD  NC51 clk n141 n51 n13 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_5_ VSS VDD  NC50 clk n141 n54 n12 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_4_ VSS VDD  NC49 clk n141 n74 n11 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_3_ VSS VDD  NC48 clk n141 n68 n10 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_2_ VSS VDD  NC47 clk n141 n55 n9 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_1_ VSS VDD  NC46 clk n141 n50 n8 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_0_ VSS VDD  NC45 clk n141 n64 n7 ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg VSS VDD  n136 clk n141 n43 n5 ASYNC_DFFHx1_ASAP7_75t_R
Xmult_x_4_U39 VSS VDD  mult_x_4_n49 mult_x_4_n52 n94 mult_x_4_n34 mult_x_4_n35 FAx1_ASAP7_75t_R
Xmult_x_4_U35 VSS VDD  mult_x_4_n36 mult_x_4_n45 mult_x_4_n32 mult_x_4_n29 mult_x_4_n30 FAx1_ASAP7_75t_R
Xmult_x_4_U32 VSS VDD  mult_x_4_n41 mult_x_4_n44 mult_x_4_n31 mult_x_4_n25 mult_x_4_n26 FAx1_ASAP7_75t_R
XU61 VSS VDD  n138 n88 INVx3_ASAP7_75t_R
XU62 VSS VDD  n86 n139 INVx3_ASAP7_75t_R
XU63 VSS VDD  n82 n44 INVx2_ASAP7_75t_R
XU64 VSS VDD  n79 n122 INVx2_ASAP7_75t_R
XU65 VSS VDD  n32 n37 mult_x_4_n49 NOR2x2_ASAP7_75t_R
XU66 VSS VDD  n38 n31 mult_x_4_n52 NOR2x1_ASAP7_75t_R
XU67 VSS VDD  n32 n36 n31 n37 n94 NOR4xp75_ASAP7_75t_R
XU68 VSS VDD  n88 n139 n136 AND2x6_ASAP7_75t_R
XU69 VSS VDD  n24 n79 BUFx5_ASAP7_75t_R
XU70 VSS VDD  mult_x_4_n35 n82 BUFx4_ASAP7_75t_R
XU71 VSS VDD  n34 n38 n32 n36 mult_x_4_n31 NOR4xp75_ASAP7_75t_R
XU72 VSS VDD  n34 n37 mult_x_4_n41 NOR2x1_ASAP7_75t_R
XU73 VSS VDD  mult_x_4_n25 n48 INVx1_ASAP7_75t_R
XU74 VSS VDD  n39 n138 BUFx5_ASAP7_75t_R
XU75 VSS VDD  n40 n86 BUFx5_ASAP7_75t_R
XU76 VSS VDD  n38 n33 mult_x_4_n44 NOR2x1_ASAP7_75t_R
XU77 VSS VDD  n81 n128 INVx2_ASAP7_75t_R
XU78 VSS VDD  n77 n132 INVx2_ASAP7_75t_R
XU79 VSS VDD  n47 TIEHIx1_ASAP7_75t_R
XU80 VSS VDD  n47 out[8] INVxp33_ASAP7_75t_R
XU81 VSS VDD  n47 out[9] INVxp33_ASAP7_75t_R
XU82 VSS VDD  n93 n105 n106 NOR2xp33_ASAP7_75t_R
XU83 VSS VDD  n136 n95 INVx5_ASAP7_75t_R
XU84 VSS VDD  rst_n n49 INVx8_ASAP7_75t_R
XU85 VSS VDD  rst_n n50 INVx8_ASAP7_75t_R
XU86 VSS VDD  rst_n n51 INVx8_ASAP7_75t_R
XU87 VSS VDD  rst_n n52 INVx8_ASAP7_75t_R
XU88 VSS VDD  rst_n n53 INVx8_ASAP7_75t_R
XU89 VSS VDD  rst_n n54 INVx8_ASAP7_75t_R
XU90 VSS VDD  rst_n n55 INVx8_ASAP7_75t_R
XU91 VSS VDD  rst_n n56 INVx8_ASAP7_75t_R
XU92 VSS VDD  rst_n n57 INVx8_ASAP7_75t_R
XU93 VSS VDD  rst_n n58 INVx8_ASAP7_75t_R
XU94 VSS VDD  rst_n n59 INVx8_ASAP7_75t_R
XU95 VSS VDD  rst_n n60 INVx8_ASAP7_75t_R
XU96 VSS VDD  rst_n n61 INVx8_ASAP7_75t_R
XU97 VSS VDD  rst_n n62 INVx8_ASAP7_75t_R
XU98 VSS VDD  rst_n n63 INVx8_ASAP7_75t_R
XU99 VSS VDD  rst_n n64 INVx8_ASAP7_75t_R
XU100 VSS VDD  rst_n n65 INVx8_ASAP7_75t_R
XU101 VSS VDD  rst_n n66 INVx8_ASAP7_75t_R
XU102 VSS VDD  rst_n n67 INVx8_ASAP7_75t_R
XU103 VSS VDD  rst_n n68 INVx8_ASAP7_75t_R
XU104 VSS VDD  rst_n n69 INVx8_ASAP7_75t_R
XU105 VSS VDD  n107 n106 n76 OR2x2_ASAP7_75t_R
XU106 VSS VDD  rst_n n70 INVx8_ASAP7_75t_R
XU107 VSS VDD  rst_n n71 INVx8_ASAP7_75t_R
XU108 VSS VDD  rst_n n72 INVx8_ASAP7_75t_R
XU109 VSS VDD  rst_n n73 INVx8_ASAP7_75t_R
XU110 VSS VDD  n123 n90 INVx4_ASAP7_75t_R
XU111 VSS VDD  n16 n123 BUFx5_ASAP7_75t_R
XU112 VSS VDD  n134 n87 INVx3_ASAP7_75t_R
XU113 VSS VDD  rst_n n74 INVx8_ASAP7_75t_R
XU114 VSS VDD  rst_n n75 INVx8_ASAP7_75t_R
XU115 VSS VDD  n107 n106 n113 NOR2xp33_ASAP7_75t_R
XU116 VSS VDD  n20 n77 BUFx5_ASAP7_75t_R
XU117 VSS VDD  rst_n n78 INVx8_ASAP7_75t_R
XU118 VSS VDD  rst_n n80 INVx8_ASAP7_75t_R
XU119 VSS VDD  n18 n81 BUFx5_ASAP7_75t_R
XU120 VSS VDD  rst_n n83 INVx8_ASAP7_75t_R
XU121 VSS VDD  rst_n n84 INVx8_ASAP7_75t_R
XU122 VSS VDD  rst_n n85 INVx8_ASAP7_75t_R
XU123 VSS VDD  n30 n134 BUFx5_ASAP7_75t_R
XU124 VSS VDD  mult_x_4_n41 mult_x_4_n44 mult_x_4_n31 n89 MAJIxp5_ASAP7_75t_R
XU125 VSS VDD  n28 n131 BUFx5_ASAP7_75t_R
XU126 VSS VDD  n131 n91 INVx4_ASAP7_75t_R
XU127 VSS VDD  n26 n127 BUFx5_ASAP7_75t_R
XU128 VSS VDD  n127 n92 INVx4_ASAP7_75t_R
XU129 VSS VDD  n32 n36 n31 n37 n93 NOR4xp25_ASAP7_75t_R
XU130 VSS VDD  n32 n36 n31 n37 mult_x_4_n38 OR4x2_ASAP7_75t_R
XU131 VSS VDD  rst_n n96 INVx8_ASAP7_75t_R
XU132 VSS VDD  rst_n n97 INVx8_ASAP7_75t_R
XU133 VSS VDD  rst_n n43 INVx8_ASAP7_75t_R
XU134 VSS VDD  n141 TIELOx1_ASAP7_75t_R
XU135 VSS VDD  n7 out[0] INVxp33_ASAP7_75t_R
XU136 VSS VDD  n9 out[2] INVxp33_ASAP7_75t_R
XU137 VSS VDD  n8 out[1] INVxp33_ASAP7_75t_R
XU138 VSS VDD  n5 out_valid INVxp33_ASAP7_75t_R
XU139 VSS VDD  n12 out[5] INVxp33_ASAP7_75t_R
XU140 VSS VDD  n13 out[6] INVxp33_ASAP7_75t_R
XU141 VSS VDD  n14 out[7] INVxp33_ASAP7_75t_R
XU142 VSS VDD  n10 out[3] INVxp33_ASAP7_75t_R
XU143 VSS VDD  n11 out[4] INVxp33_ASAP7_75t_R
XU144 VSS VDD  n38 n32 n99 NOR2xp33_ASAP7_75t_R
XU145 VSS VDD  n34 n36 n98 NOR2xp33_ASAP7_75t_R
XU146 VSS VDD  n99 n98 n100 NOR2xp33_ASAP7_75t_R
XU147 VSS VDD  mult_x_4_n31 n100 mult_x_4_n32 NOR2xp33_ASAP7_75t_R
XU148 VSS VDD  n34 n36 n35 n33 mult_x_4_n36 NOR4xp25_ASAP7_75t_R
XU149 VSS VDD  n37 n33 mult_x_4_n45 NOR2xp33_ASAP7_75t_R
XU150 VSS VDD  n31 n35 NC28 NOR2xp33_ASAP7_75t_R
XU151 VSS VDD  n36 n31 n102 NOR2xp33_ASAP7_75t_R
XU152 VSS VDD  n32 n35 n101 NOR2xp33_ASAP7_75t_R
XU153 VSS VDD  n102 n101 NC29 XOR2xp5_ASAP7_75t_R
XU154 VSS VDD  n35 n33 n109 NOR2xp33_ASAP7_75t_R
XU155 VSS VDD  n32 n36 n104 NOR2xp33_ASAP7_75t_R
XU156 VSS VDD  NC28 n104 mult_x_4_n38 n115 NAND3xp33_ASAP7_75t_R
XU157 VSS VDD  n35 n32 n36 n107 NOR3xp33_ASAP7_75t_R
XU158 VSS VDD  n31 n37 n103 NOR2xp33_ASAP7_75t_R
XU159 VSS VDD  n104 n103 n105 NOR2xp33_ASAP7_75t_R
XU160 VSS VDD  n76 n115 n108 NAND2xp33_ASAP7_75t_R
XU161 VSS VDD  n109 n108 A0  NC30 HAxp5_ASAP7_75t_R
XU162 VSS VDD  n36 n33 n111 NOR2xp33_ASAP7_75t_R
XU163 VSS VDD  n34 n35 n110 NOR2xp33_ASAP7_75t_R
XU164 VSS VDD  n111 n110 n112 NOR2xp33_ASAP7_75t_R
XU165 VSS VDD  mult_x_4_n36 n112 n117 NOR2xp33_ASAP7_75t_R
XU166 VSS VDD  n33 n35 n113 n114 OR3x1_ASAP7_75t_R
XU167 VSS VDD  n115 n114 n116 NAND2xp33_ASAP7_75t_R
XU168 VSS VDD  n116 n117 n82 A1  NC31 FAx1_ASAP7_75t_R
XU169 VSS VDD  n44 n116 n117 n118 MAJIxp5_ASAP7_75t_R
XU170 VSS VDD  mult_x_4_n30 n118 mult_x_4_n34 A2  NC32 FAx1_ASAP7_75t_R
XU171 VSS VDD  mult_x_4_n30 n118 mult_x_4_n34 n119 MAJx2_ASAP7_75t_R
XU172 VSS VDD  mult_x_4_n29 n119 mult_x_4_n26 A3  NC33 FAx1_ASAP7_75t_R
XU173 VSS VDD  n34 n38 n121 NOR2xp33_ASAP7_75t_R
XU174 VSS VDD  mult_x_4_n29 n119 mult_x_4_n26 n120 MAJIxp5_ASAP7_75t_R
XU175 VSS VDD  n89 n121 n120 A4  NC34 FAx1_ASAP7_75t_R
XU176 VSS VDD  n48 n121 n120 NC35 MAJx2_ASAP7_75t_R
XU177 VSS VDD  n23 n15 NC36 XOR2xp5_ASAP7_75t_R
XU178 VSS VDD  n23 n15 n124 NOR2xp33_ASAP7_75t_R
XU179 VSS VDD  n79 n124 n90 A5  NC37 FAx1_ASAP7_75t_R
XU180 VSS VDD  n90 n124 n122 n125 MAJIxp5_ASAP7_75t_R
XU181 VSS VDD  n17 n25 n125 A6  NC38 FAx1_ASAP7_75t_R
XU182 VSS VDD  n17 n25 n125 n126 MAJIxp5_ASAP7_75t_R
XU183 VSS VDD  n81 n126 n92 A7  NC39 FAx1_ASAP7_75t_R
XU184 VSS VDD  n128 n126 n92 n129 MAJIxp5_ASAP7_75t_R
XU185 VSS VDD  n19 n27 n129 A8  NC40 FAx1_ASAP7_75t_R
XU186 VSS VDD  n19 n27 n129 n130 MAJIxp5_ASAP7_75t_R
XU187 VSS VDD  n77 n130 n91 A9  NC41 FAx1_ASAP7_75t_R
XU188 VSS VDD  n132 n130 n91 n133 MAJIxp5_ASAP7_75t_R
XU189 VSS VDD  n29 n133 n21 A10  NC42 FAx1_ASAP7_75t_R
XU190 VSS VDD  n29 n133 n21 n135 MAJIxp5_ASAP7_75t_R
XU191 VSS VDD  n135 n22 n87 A11  NC43 FAx1_ASAP7_75t_R
XU192 VSS VDD  in_valid in1_IFM[0] NC18 AND2x2_ASAP7_75t_R
XU193 VSS VDD  in_valid in1_IFM[1] NC19 AND2x2_ASAP7_75t_R
XU194 VSS VDD  in_valid in1_IFM[2] NC20 AND2x2_ASAP7_75t_R
XU195 VSS VDD  in_valid in1_IFM[3] NC21 AND2x2_ASAP7_75t_R
XU196 VSS VDD  in_valid in2_IFM[0] NC22 AND2x2_ASAP7_75t_R
XU197 VSS VDD  in_valid in2_IFM[1] NC23 AND2x2_ASAP7_75t_R
XU198 VSS VDD  in_valid in2_IFM[2] NC24 AND2x2_ASAP7_75t_R
XU199 VSS VDD  in_valid in2_IFM[3] NC25 AND2x2_ASAP7_75t_R
XU200 VSS VDD  n95 n23 NC45 NOR2xp33_ASAP7_75t_R
XU201 VSS VDD  n95 n79 NC46 NOR2xp33_ASAP7_75t_R
XU202 VSS VDD  n95 n25 NC47 NOR2xp33_ASAP7_75t_R
XU203 VSS VDD  n127 n95 NC48 NOR2xp33_ASAP7_75t_R
XU204 VSS VDD  n95 n27 NC49 NOR2xp33_ASAP7_75t_R
XU205 VSS VDD  n131 n95 NC50 NOR2xp33_ASAP7_75t_R
XU206 VSS VDD  n95 n29 NC51 NOR2xp33_ASAP7_75t_R
XU207 VSS VDD  n134 n95 NC52 NOR2xp33_ASAP7_75t_R
XU208 VSS VDD  n88 in_valid n137 NOR2xp33_ASAP7_75t_R
XU209 VSS VDD  n139 n137 n42 NOR2xp33_ASAP7_75t_R
XU210 VSS VDD  n139 n88 n140 NOR2xp33_ASAP7_75t_R
XU211 VSS VDD  n136 n140 n41 NOR2xp33_ASAP7_75t_R
.ENDS