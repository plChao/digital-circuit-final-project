.SUBCKT MAC VSS VDD  in1_IFM[3] in1_IFM[2] in1_IFM[1] in1_IFM[0] in2_IFM[3] in2_IFM[2] in2_IFM[1] in2_IFM[0] out[9] out[8] out[7] out[6] out[5] out[4] out[3] out[2] out[1] out[0] clk rst_n in_valid out_valid
Xcstate_reg_0_ VSS VDD  n108 clk n238 n138 n106 ASYNC_DFFHx1_ASAP7_75t_R
Xcstate_reg_1_ VSS VDD  n107 clk n238 n128 n105 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_3_ VSS VDD  N25 clk n238 n167 n104 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_2_ VSS VDD  N24 clk n238 n148 n103 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_1_ VSS VDD  N23 clk n238 n125 n102 ASYNC_DFFHx1_ASAP7_75t_R
Xin2_reg_0_ VSS VDD  N22 clk n238 n119 n101 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_3_ VSS VDD  N21 clk n238 n124 n100 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_2_ VSS VDD  N20 clk n238 n121 n99 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_1_ VSS VDD  N19 clk n238 n116 n98 ASYNC_DFFHx1_ASAP7_75t_R
Xin1_reg_0_ VSS VDD  N18 clk n238 n156 n97 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_7_ VSS VDD  add_x_7_n6 clk n238 n145 n96 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_6_ VSS VDD  add_x_8_n6 clk n238 n137 n95 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_5_ VSS VDD  add_x_9_n6 clk n238 n154 n94 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_4_ VSS VDD  add_x_10_n6 clk n238 n146 n93 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_3_ VSS VDD  add_x_11_n6 clk n238 n142 n92 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_2_ VSS VDD  add_x_12_n6 clk n238 n122 n91 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_1_ VSS VDD  add_x_6_n6 clk n238 n141 n90 ASYNC_DFFHx1_ASAP7_75t_R
Xfprod_1_reg_0_ VSS VDD  fprod_0_ clk n238 n131 n89 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_8_ VSS VDD  temp_1 clk n238 n117 n88 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_7_ VSS VDD  temp_0[7] clk n238 n129 n87 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_6_ VSS VDD  temp_0[6] clk n238 n140 n86 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_5_ VSS VDD  temp_0[5] clk n238 n157 n85 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_4_ VSS VDD  temp_0[4] clk n238 n127 n84 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_3_ VSS VDD  temp_0[3] clk n238 n126 n83 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_2_ VSS VDD  temp_0[2] clk n238 n155 n82 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_1_ VSS VDD  temp_0[1] clk n238 n115 n81 ASYNC_DFFHx1_ASAP7_75t_R
Xsum_reg_0_ VSS VDD  temp_0[0] clk n238 n166 n80 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_8_ VSS VDD  N37 clk n238 n130 n79 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_7_ VSS VDD  N36 clk n238 n151 n78 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_6_ VSS VDD  N35 clk n238 n123 n77 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_5_ VSS VDD  N34 clk n238 n118 n76 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_4_ VSS VDD  N33 clk n238 n120 n75 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_3_ VSS VDD  N32 clk n238 n147 n74 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_2_ VSS VDD  N31 clk n238 n144 n73 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_1_ VSS VDD  N30 clk n238 n132 n72 ASYNC_DFFHx1_ASAP7_75t_R
Xout_reg_0_ VSS VDD  N29 clk n238 n139 n71 ASYNC_DFFHx1_ASAP7_75t_R
Xout_valid_reg VSS VDD  n218 clk n238 n109 n69 ASYNC_DFFHx1_ASAP7_75t_R
XU128 VSS VDD  n143 n226 add_x_9_n6 NOR2xp33_ASAP7_75t_R
XU129 VSS VDD  in_valid in2_IFM[1] N23 AND2x2_ASAP7_75t_R
XU130 VSS VDD  in_valid in2_IFM[2] N24 AND2x2_ASAP7_75t_R
XU131 VSS VDD  in_valid in2_IFM[0] N22 AND2x2_ASAP7_75t_R
XU132 VSS VDD  in_valid in2_IFM[3] N25 AND2x2_ASAP7_75t_R
XU133 VSS VDD  in_valid in1_IFM[2] N20 AND2x2_ASAP7_75t_R
XU134 VSS VDD  in_valid in1_IFM[1] N19 AND2x2_ASAP7_75t_R
XU135 VSS VDD  in_valid in1_IFM[0] N18 AND2x2_ASAP7_75t_R
XU136 VSS VDD  n235 n162 INVx3_ASAP7_75t_R
XU137 VSS VDD  n158 n236 INVx3_ASAP7_75t_R
XU138 VSS VDD  n195 n194 n223 NOR2xp33_ASAP7_75t_R
XU139 VSS VDD  n134 n183 n188 NOR2xp33_ASAP7_75t_R
XU140 VSS VDD  n104 n99 n189 NOR2xp33_ASAP7_75t_R
XU141 VSS VDD  n100 n103 n190 NOR2xp33_ASAP7_75t_R
XU142 VSS VDD  n181 n180 n159 XOR2xp5_ASAP7_75t_R
XU143 VSS VDD  n173 n172 n191 NOR2xp33_ASAP7_75t_R
XU144 VSS VDD  n111 TIEHIx1_ASAP7_75t_R
XU145 VSS VDD  n111 out[9] INVx1_ASAP7_75t_R
XU146 VSS VDD  n218 n112 INVx4_ASAP7_75t_R
XU147 VSS VDD  n162 n236 n218 AND2x6_ASAP7_75t_R
XU148 VSS VDD  n105 n235 BUFx5_ASAP7_75t_R
XU149 VSS VDD  n106 n158 BUFx5_ASAP7_75t_R
XU150 VSS VDD  n186 n185 n187 NOR2xp33_ASAP7_75t_R
XU151 VSS VDD  n103 n98 n177 NOR2xp33_ASAP7_75t_R
XU152 VSS VDD  n202 n201 n227 NOR2xp33_ASAP7_75t_R
XU153 VSS VDD  in_valid in1_IFM[3] N21 AND2x2_ASAP7_75t_R
XU154 VSS VDD  n150 n203 add_x_7_n6 NAND2xp5_ASAP7_75t_R
XU155 VSS VDD  n233 n219 n221 NAND2xp5_ASAP7_75t_R
XU156 VSS VDD  n152 n207 INVx2_ASAP7_75t_R
XU157 VSS VDD  n190 n189 n161 NAND2xp5_ASAP7_75t_R
XU158 VSS VDD  n149 n215 INVx2_ASAP7_75t_R
XU159 VSS VDD  n153 n211 INVx2_ASAP7_75t_R
XU160 VSS VDD  n181 n180 n160 XNOR2xp5_ASAP7_75t_R
XU161 VSS VDD  n188 n187 n199 XNOR2xp5_ASAP7_75t_R
XU162 VSS VDD  n179 n184 n113 XOR2xp5_ASAP7_75t_R
XU163 VSS VDD  n179 n184 n197 XNOR2xp5_ASAP7_75t_R
XU164 VSS VDD  n225 n224 n114 NAND2xp33_ASAP7_75t_R
XU165 VSS VDD  rst_n n115 INVx8_ASAP7_75t_R
XU166 VSS VDD  rst_n n116 INVx8_ASAP7_75t_R
XU167 VSS VDD  rst_n n117 INVx8_ASAP7_75t_R
XU168 VSS VDD  rst_n n118 INVx8_ASAP7_75t_R
XU169 VSS VDD  rst_n n119 INVx8_ASAP7_75t_R
XU170 VSS VDD  rst_n n120 INVx8_ASAP7_75t_R
XU171 VSS VDD  rst_n n121 INVx8_ASAP7_75t_R
XU172 VSS VDD  rst_n n122 INVx8_ASAP7_75t_R
XU173 VSS VDD  rst_n n123 INVx8_ASAP7_75t_R
XU174 VSS VDD  rst_n n124 INVx8_ASAP7_75t_R
XU175 VSS VDD  rst_n n125 INVx8_ASAP7_75t_R
XU176 VSS VDD  rst_n n126 INVx8_ASAP7_75t_R
XU177 VSS VDD  rst_n n127 INVx8_ASAP7_75t_R
XU178 VSS VDD  rst_n n128 INVx8_ASAP7_75t_R
XU179 VSS VDD  rst_n n129 INVx8_ASAP7_75t_R
XU180 VSS VDD  rst_n n130 INVx8_ASAP7_75t_R
XU181 VSS VDD  rst_n n131 INVx8_ASAP7_75t_R
XU182 VSS VDD  rst_n n132 INVx8_ASAP7_75t_R
XU183 VSS VDD  n188 n187 n133 XOR2xp5_ASAP7_75t_R
XU184 VSS VDD  n221 n220 n134 NOR2xp33_ASAP7_75t_R
XU185 VSS VDD  n182 n159 n135 XOR2xp5_ASAP7_75t_R
XU186 VSS VDD  n225 n224 n143 AND2x2_ASAP7_75t_R
XU187 VSS VDD  n190 n189 n136 AND2x2_ASAP7_75t_R
XU188 VSS VDD  rst_n n137 INVx8_ASAP7_75t_R
XU189 VSS VDD  rst_n n138 INVx8_ASAP7_75t_R
XU190 VSS VDD  rst_n n139 INVx8_ASAP7_75t_R
XU191 VSS VDD  rst_n n140 INVx8_ASAP7_75t_R
XU192 VSS VDD  rst_n n141 INVx8_ASAP7_75t_R
XU193 VSS VDD  rst_n n142 INVx8_ASAP7_75t_R
XU194 VSS VDD  n188 n161 n150 OR2x2_ASAP7_75t_R
XU195 VSS VDD  rst_n n144 INVx8_ASAP7_75t_R
XU196 VSS VDD  rst_n n145 INVx8_ASAP7_75t_R
XU197 VSS VDD  n221 n220 n184 OR2x2_ASAP7_75t_R
XU198 VSS VDD  n182 n159 n196 XNOR2xp5_ASAP7_75t_R
XU199 VSS VDD  rst_n n146 INVx8_ASAP7_75t_R
XU200 VSS VDD  rst_n n147 INVx8_ASAP7_75t_R
XU201 VSS VDD  rst_n n148 INVx8_ASAP7_75t_R
XU202 VSS VDD  n95 n149 BUFx5_ASAP7_75t_R
XU203 VSS VDD  rst_n n151 INVx8_ASAP7_75t_R
XU204 VSS VDD  n91 n152 BUFx5_ASAP7_75t_R
XU205 VSS VDD  n93 n153 BUFx5_ASAP7_75t_R
XU206 VSS VDD  rst_n n154 INVx8_ASAP7_75t_R
XU207 VSS VDD  rst_n n155 INVx8_ASAP7_75t_R
XU208 VSS VDD  rst_n n156 INVx8_ASAP7_75t_R
XU209 VSS VDD  rst_n n157 INVx8_ASAP7_75t_R
XU210 VSS VDD  n86 n214 BUFx5_ASAP7_75t_R
XU211 VSS VDD  n214 n163 INVx4_ASAP7_75t_R
XU212 VSS VDD  n84 n210 BUFx5_ASAP7_75t_R
XU213 VSS VDD  n210 n164 INVx4_ASAP7_75t_R
XU214 VSS VDD  n82 n206 BUFx5_ASAP7_75t_R
XU215 VSS VDD  n206 n165 INVx4_ASAP7_75t_R
XU216 VSS VDD  rst_n n166 INVx8_ASAP7_75t_R
XU217 VSS VDD  rst_n n167 INVx8_ASAP7_75t_R
XU218 VSS VDD  rst_n n109 INVx8_ASAP7_75t_R
XU219 VSS VDD  n238 TIELOx1_ASAP7_75t_R
XU220 VSS VDD  n102 n98 n97 n101 n233 NOR4xp25_ASAP7_75t_R
XU221 VSS VDD  n103 n97 n170 NOR2xp33_ASAP7_75t_R
XU222 VSS VDD  n102 n98 n169 NOR2xp33_ASAP7_75t_R
XU223 VSS VDD  n99 n101 n168 NOR2xp33_ASAP7_75t_R
XU224 VSS VDD  n169 n168 A0  n171 HAxp5_ASAP7_75t_R
XU225 VSS VDD  n170 n171 A1  n219 HAxp5_ASAP7_75t_R
XU226 VSS VDD  n99 n102 n98 n101 n173 NOR4xp25_ASAP7_75t_R
XU227 VSS VDD  n103 n97 n171 n172 NOR3xp33_ASAP7_75t_R
XU228 VSS VDD  n104 n97 n174 NOR2xp33_ASAP7_75t_R
XU229 VSS VDD  n191 n174 A2  n193 HAxp5_ASAP7_75t_R
XU230 VSS VDD  n99 n102 n178 NOR2xp33_ASAP7_75t_R
XU231 VSS VDD  n100 n101 n176 NOR2xp33_ASAP7_75t_R
XU232 VSS VDD  n178 n176 A3  n175 HAxp5_ASAP7_75t_R
XU233 VSS VDD  n177 n175 A4  n192 HAxp5_ASAP7_75t_R
XU234 VSS VDD  n193 n192 A5  n220 HAxp5_ASAP7_75t_R
XU235 VSS VDD  n178 n177 n176 n179 MAJIxp5_ASAP7_75t_R
XU236 VSS VDD  n104 n98 n182 NOR2xp33_ASAP7_75t_R
XU237 VSS VDD  n103 n99 n181 NOR2xp33_ASAP7_75t_R
XU238 VSS VDD  n100 n102 n180 NOR2xp33_ASAP7_75t_R
XU239 VSS VDD  n197 n196 n183 NOR2xp33_ASAP7_75t_R
XU240 VSS VDD  n188 n161 n202 NOR2xp33_ASAP7_75t_R
XU241 VSS VDD  n100 n104 n228 NOR2xp33_ASAP7_75t_R
XU242 VSS VDD  n100 n103 n99 n102 n186 NOR4xp25_ASAP7_75t_R
XU243 VSS VDD  n104 n98 n160 n185 NOR3xp33_ASAP7_75t_R
XU244 VSS VDD  n190 n189 A6  n198 HAxp5_ASAP7_75t_R
XU245 VSS VDD  n198 n133 A7  n225 HAxp5_ASAP7_75t_R
XU246 VSS VDD  n104 n97 n191 n195 NOR3xp33_ASAP7_75t_R
XU247 VSS VDD  n193 n192 n194 AND2x2_ASAP7_75t_R
XU248 VSS VDD  n135 n113 A8  n222 HAxp5_ASAP7_75t_R
XU249 VSS VDD  n223 n222 n224 NOR2xp33_ASAP7_75t_R
XU250 VSS VDD  n199 n198 n200 NOR2xp33_ASAP7_75t_R
XU251 VSS VDD  n136 n200 n201 NOR2xp33_ASAP7_75t_R
XU252 VSS VDD  n143 n228 n227 n203 MAJIxp5_ASAP7_75t_R
XU253 VSS VDD  n69 out_valid INVxp33_ASAP7_75t_R
XU254 VSS VDD  n71 out[0] INVxp33_ASAP7_75t_R
XU255 VSS VDD  n73 out[2] INVxp33_ASAP7_75t_R
XU256 VSS VDD  n74 out[3] INVxp33_ASAP7_75t_R
XU257 VSS VDD  n75 out[4] INVxp33_ASAP7_75t_R
XU258 VSS VDD  n76 out[5] INVxp33_ASAP7_75t_R
XU259 VSS VDD  n77 out[6] INVxp33_ASAP7_75t_R
XU260 VSS VDD  n78 out[7] INVxp33_ASAP7_75t_R
XU261 VSS VDD  n79 out[8] INVxp33_ASAP7_75t_R
XU262 VSS VDD  n72 out[1] INVxp33_ASAP7_75t_R
XU263 VSS VDD  n80 n89 temp_0[0] XOR2xp5_ASAP7_75t_R
XU264 VSS VDD  n80 n89 n204 OR2x2_ASAP7_75t_R
XU265 VSS VDD  n81 n90 n204 A9  temp_0[1] FAx1_ASAP7_75t_R
XU266 VSS VDD  n90 n81 n204 n205 MAJIxp5_ASAP7_75t_R
XU267 VSS VDD  n152 n205 n165 A10  temp_0[2] FAx1_ASAP7_75t_R
XU268 VSS VDD  n207 n205 n165 n208 MAJIxp5_ASAP7_75t_R
XU269 VSS VDD  n92 n83 n208 A11  temp_0[3] FAx1_ASAP7_75t_R
XU270 VSS VDD  n92 n83 n208 n209 MAJIxp5_ASAP7_75t_R
XU271 VSS VDD  n153 n209 n164 A12  temp_0[4] FAx1_ASAP7_75t_R
XU272 VSS VDD  n211 n209 n164 n212 MAJIxp5_ASAP7_75t_R
XU273 VSS VDD  n94 n85 n212 A13  temp_0[5] FAx1_ASAP7_75t_R
XU274 VSS VDD  n94 n85 n212 n213 MAJIxp5_ASAP7_75t_R
XU275 VSS VDD  n149 n213 n163 A14  temp_0[6] FAx1_ASAP7_75t_R
XU276 VSS VDD  n215 n213 n163 n216 MAJIxp5_ASAP7_75t_R
XU277 VSS VDD  n87 n216 n96 A15  temp_0[7] FAx1_ASAP7_75t_R
XU278 VSS VDD  n87 n216 n96 n217 MAJIxp5_ASAP7_75t_R
XU279 VSS VDD  n88 n217 A16  temp_1 HAxp5_ASAP7_75t_R
XU280 VSS VDD  n97 n101 fprod_0_ NOR2xp33_ASAP7_75t_R
XU281 VSS VDD  n112 n80 N29 NOR2xp33_ASAP7_75t_R
XU282 VSS VDD  n112 n81 N30 NOR2xp33_ASAP7_75t_R
XU283 VSS VDD  n206 n112 N31 NOR2xp33_ASAP7_75t_R
XU284 VSS VDD  n112 n83 N32 NOR2xp33_ASAP7_75t_R
XU285 VSS VDD  n210 n112 N33 NOR2xp33_ASAP7_75t_R
XU286 VSS VDD  n112 n85 N34 NOR2xp33_ASAP7_75t_R
XU287 VSS VDD  n214 n112 N35 NOR2xp33_ASAP7_75t_R
XU288 VSS VDD  n112 n87 N36 NOR2xp33_ASAP7_75t_R
XU289 VSS VDD  n112 n88 N37 NOR2xp33_ASAP7_75t_R
XU290 VSS VDD  n233 n219 add_x_12_n6 XOR2xp5_ASAP7_75t_R
XU291 VSS VDD  n221 n220 add_x_11_n6 XOR2xp5_ASAP7_75t_R
XU292 VSS VDD  n223 n222 add_x_10_n6 XOR2xp5_ASAP7_75t_R
XU293 VSS VDD  n225 n224 n226 NOR2xp33_ASAP7_75t_R
XU294 VSS VDD  n228 n227 n229 XOR2xp5_ASAP7_75t_R
XU295 VSS VDD  n229 n114 A17  add_x_8_n6 HAxp5_ASAP7_75t_R
XU296 VSS VDD  n98 n101 n231 NOR2xp33_ASAP7_75t_R
XU297 VSS VDD  n102 n97 n230 NOR2xp33_ASAP7_75t_R
XU298 VSS VDD  n231 n230 n232 NOR2xp33_ASAP7_75t_R
XU299 VSS VDD  n233 n232 add_x_6_n6 NOR2xp33_ASAP7_75t_R
XU300 VSS VDD  n162 in_valid n234 NOR2xp33_ASAP7_75t_R
XU301 VSS VDD  n236 n234 n108 NOR2xp33_ASAP7_75t_R
XU302 VSS VDD  n236 n162 n237 NOR2xp33_ASAP7_75t_R
XU303 VSS VDD  n218 n237 n107 NOR2xp33_ASAP7_75t_R
.ENDS


